library ieee;
use ieee.std_logic_1164.all;

package register_file_types is

  type reg_array is (natural range <>) of std_logic_vector;

end package;
