library ieee;
use ieee.std_logic_1164.all;

use work.my_arith_functions.all;

package p4_carries_logic_network_types is

end package;
